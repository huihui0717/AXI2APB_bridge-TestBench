`ifndef X2P_ENV__SV
`define X2P_ENV__SV

class x2p_env extends uvm_env;






endclass: x2p_env

`endif  // X2P_ENV__SV
