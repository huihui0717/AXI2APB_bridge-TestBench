module test;





endmodule
