module top();







endmodule: top
