`ifndef  AXI_PACKET__SV
`define  AXI_PACKET__SV

class axi_packet;





endclass: axi_packet





`endif  // AXI_PACKET__SV
